library ieee; 
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.globals.all;

entity P4_ADDER is
    port ( 
        A : in std_logic_vector(WORD_SIZE_c-1 downto 0);
        B : in std_logic_vector(WORD_SIZE_c-1 downto 0);
        C_in : in std_logic;
        S: out std_logic_vector(WORD_SIZE_c-1 downto 0);
        C_out : out std_logic
    );
end P4_ADDER;

architecture STRUCTURAL of P4_ADDER is

    --------------------------------------------------
    -- Component declarations
    --------------------------------------------------

    -- Carry generator circuit
    component CARRY_GENERATOR_GEN is
        generic(
            NBIT_IN : integer; -- Number of bits of input
            NCARRY : integer; -- Number of carries generated by this block
            NBIT_CARRY : integer -- Number of bits for a carry
        );
        port (
            A : in std_logic_vector(NBIT_IN-1 downto 0);
            B : in std_logic_vector(NBIT_IN-1 downto 0);
            C_in : in std_logic;
            O : out std_logic_vector(NCARRY-1 downto 0)
        ) ;
    end component ;

    -- Generic 2to1 multiplexer
    component MUX21_GEN is
        generic (NBIT: integer);
        port (A: in std_logic_vector(NBIT-1 downto 0) ;
              B: in std_logic_vector(NBIT-1 downto 0);
              SEL: in std_logic;
              Y: out std_logic_vector(NBIT-1 downto 0));
    end component;

    -- Generic RCA
    component RCA_GEN is 
        generic(NBIT: integer);
        port (A: in std_logic_vector(NBIT-1 downto 0);
              B: in std_logic_vector(NBIT-1 downto 0);
              C_in: in std_logic;
              S: out std_logic_vector(NBIT-1 downto 0);
              C_out: out std_logic);
    end component;

    --------------------------------------------------
    -- Signals declarations
    --------------------------------------------------
    type S_PART_t is array(ADDER_CARRY_NUMBER_c-1 downto 0) of std_logic_vector(ADDER_CARRY_SIZE_c-1 downto 0);
    signal S_C_IN_0 : S_PART_t;
    signal S_C_IN_1 : S_PART_t;
    signal C_SEL_i : std_logic_vector(ADDER_CARRY_NUMBER_c-1 downto 0);

begin

    CARRY_GENERATOR_GEN_I : CARRY_GENERATOR_GEN
    generic map(
        NBIT_IN => WORD_SIZE_c,
        NCARRY => ADDER_CARRY_NUMBER_c,
        NBIT_CARRY => ADDER_CARRY_SIZE_c
    )
    port map(
        A => A,
        B => B,
        C_in => C_in,
        O => C_SEL_i
    );

    RCA_FIRST : RCA_GEN
    generic map (
        NBIT => ADDER_CARRY_SIZE_c)
    port map (
        A => A(ADDER_CARRY_SIZE_c-1 downto 0),
        B => B(ADDER_CARRY_SIZE_c-1 downto 0),
        C_in => C_in,
        S => S(ADDER_CARRY_SIZE_c-1 downto 0),
        C_out => open);

    ADDER_I : for I in 1 to ADDER_CARRY_NUMBER_c-1 generate

        -- '0' carry in RCA
        RCA_GEN_0 : RCA_GEN
        generic map (
            NBIT => ADDER_CARRY_SIZE_c)
        port map (
            A => A((I+1)*ADDER_CARRY_SIZE_c-1 downto I*ADDER_CARRY_SIZE_c),
            B => B((I+1)*ADDER_CARRY_SIZE_c-1 downto I*ADDER_CARRY_SIZE_c),
            C_in => '0',
            S => S_C_IN_0(I),
            C_out => open);

        -- '1' carry in RCA
        RCA_GEN_1 : RCA_GEN
        generic map (
            NBIT => ADDER_CARRY_SIZE_c)
        port map (
            A => A((I+1)*ADDER_CARRY_SIZE_c-1 downto I*ADDER_CARRY_SIZE_c),
            B => B((I+1)*ADDER_CARRY_SIZE_c-1 downto I*ADDER_CARRY_SIZE_c),
            C_in => '1',
            S => S_C_IN_1(I),
            C_out => open);

        -- Select the correct result
        MUX21_GEN_0 : MUX21_GEN
        generic map (
            NBIT => ADDER_CARRY_SIZE_c)
        port map (
            A => S_C_IN_0(I),
            B => S_C_IN_1(I),
            SEL => C_SEL_i(I-1),
            Y => S((I+1)*ADDER_CARRY_SIZE_c-1 downto I*ADDER_CARRY_SIZE_c));

    end generate;


    C_out <= C_SEL_i(ADDER_CARRY_NUMBER_c-1);

end STRUCTURAL;
